`ifndef COM
`define COM

class apb_common;
  static int num_matches;
  static int num_mismatches;
  static int total_pkt_count;
endclass

`endif
